
module PG_generate_0 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module CUS_PLUS_0 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n2;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n2), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n2) );
endmodule


module Carry_Generate_0 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n2) );
endmodule


module SUM_generate_0 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module PG_generate_1 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_2 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_3 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_4 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_5 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_6 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_7 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_8 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_9 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_10 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_11 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_12 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_13 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_14 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module PG_generate_15 ( add_1, add_2, Propagate, Generate );
  input add_1, add_2;
  output Propagate, Generate;


  XOR2_X1 U2 ( .A(add_2), .B(add_1), .Z(Propagate) );
  AND2_X1 U1 ( .A1(add_2), .A2(add_1), .ZN(Generate) );
endmodule


module CUS_PLUS_1 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_2 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_3 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_4 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_5 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_6 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AOI21_X1 U1 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
  AND2_X1 U2 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U3 ( .A(n1), .ZN(alpha[0]) );
endmodule


module CUS_PLUS_7 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AOI21_X1 U1 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
  AND2_X1 U2 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U3 ( .A(n1), .ZN(alpha[0]) );
endmodule


module CUS_PLUS_8 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_9 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_10 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_11 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_12 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_13 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_14 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_15 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_16 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_17 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_18 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_19 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_20 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_21 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_22 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_23 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_24 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  AND2_X1 U1 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
  INV_X1 U2 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U3 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
endmodule


module CUS_PLUS_25 ( g_high, g_low, p_high, p_low, alpha, beta );
  input [0:0] g_high;
  input [0:0] g_low;
  input [0:0] p_high;
  input [0:0] p_low;
  output [0:0] alpha;
  output [0:0] beta;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(alpha[0]) );
  AOI21_X1 U2 ( .B1(g_low[0]), .B2(p_high[0]), .A(g_high[0]), .ZN(n1) );
  AND2_X1 U3 ( .A1(p_low[0]), .A2(p_high[0]), .ZN(beta[0]) );
endmodule


module Carry_Generate_1 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_2 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_3 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_4 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_5 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_6 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_7 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_8 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_9 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_10 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_11 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_12 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_13 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_14 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module Carry_Generate_15 ( alpha, beta, c_in, c_out );
  input [0:0] alpha;
  input [0:0] beta;
  input [0:0] c_in;
  output [0:0] c_out;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(c_out[0]) );
  AOI21_X1 U2 ( .B1(c_in[0]), .B2(beta[0]), .A(alpha[0]), .ZN(n1) );
endmodule


module SUM_generate_1 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_2 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_3 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_4 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_5 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_6 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_7 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_8 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_9 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_10 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_11 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_12 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_13 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_14 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module SUM_generate_15 ( Propagate, c_in, Sum );
  input [0:0] Propagate;
  input [0:0] c_in;
  output [0:0] Sum;


  XOR2_X1 U1 ( .A(c_in[0]), .B(Propagate[0]), .Z(Sum[0]) );
endmodule


module PPA ( add_1, add_2, c_in, sum, c_out );
  input [16:1] add_1;
  input [16:1] add_2;
  output [16:1] sum;
  output [0:0] c_out;
  input c_in;
  wire   stage_1_alpha_16_, stage_1_alpha_14, stage_1_alpha_12,
         stage_1_alpha_10, stage_1_alpha_8, stage_1_alpha_6, stage_1_alpha_4,
         stage_1_alpha_2, stage_1_beta_16_, stage_1_beta_14, stage_1_beta_12,
         stage_1_beta_10, stage_1_beta_8, stage_1_beta_6, stage_1_beta_4,
         stage_1_beta_2, stage_2_alpha_16_, stage_2_alpha_12, stage_2_alpha_8,
         stage_2_alpha_4, stage_2_beta_16_, stage_2_beta_12, stage_2_beta_8,
         stage_2_beta_4, stage_3_alpha_16_, stage_3_alpha_8, stage_3_beta_16_,
         stage_3_beta_8, stage_4_alpha_16_, stage_4_alpha_12, stage_4_beta_16_,
         stage_4_beta_12, stage_5_alpha_14_, stage_5_alpha_10, stage_5_alpha_6,
         stage_5_beta_14_, stage_5_beta_10, stage_5_beta_6, stage_6_alpha_15_,
         stage_6_alpha_13, stage_6_alpha_11, stage_6_alpha_9, stage_6_alpha_7,
         stage_6_alpha_5, stage_6_alpha_3, stage_6_beta_15_, stage_6_beta_13,
         stage_6_beta_11, stage_6_beta_9, stage_6_beta_7, stage_6_beta_5,
         stage_6_beta_3;
  wire   [15:1] Carry;
  wire   [16:1] Generate;
  wire   [16:1] Propagate;

  PG_generate_0 PG_GEN_1__PG_generate_inst ( .add_1(add_1[1]), .add_2(add_2[1]), .Propagate(Propagate[1]), .Generate(Generate[1]) );
  PG_generate_15 PG_GEN_2__PG_generate_inst ( .add_1(add_1[2]), .add_2(
        add_2[2]), .Propagate(Propagate[2]), .Generate(Generate[2]) );
  PG_generate_14 PG_GEN_3__PG_generate_inst ( .add_1(add_1[3]), .add_2(
        add_2[3]), .Propagate(Propagate[3]), .Generate(Generate[3]) );
  PG_generate_13 PG_GEN_4__PG_generate_inst ( .add_1(add_1[4]), .add_2(
        add_2[4]), .Propagate(Propagate[4]), .Generate(Generate[4]) );
  PG_generate_12 PG_GEN_5__PG_generate_inst ( .add_1(add_1[5]), .add_2(
        add_2[5]), .Propagate(Propagate[5]), .Generate(Generate[5]) );
  PG_generate_11 PG_GEN_6__PG_generate_inst ( .add_1(add_1[6]), .add_2(
        add_2[6]), .Propagate(Propagate[6]), .Generate(Generate[6]) );
  PG_generate_10 PG_GEN_7__PG_generate_inst ( .add_1(add_1[7]), .add_2(
        add_2[7]), .Propagate(Propagate[7]), .Generate(Generate[7]) );
  PG_generate_9 PG_GEN_8__PG_generate_inst ( .add_1(add_1[8]), .add_2(add_2[8]), .Propagate(Propagate[8]), .Generate(Generate[8]) );
  PG_generate_8 PG_GEN_9__PG_generate_inst ( .add_1(add_1[9]), .add_2(add_2[9]), .Propagate(Propagate[9]), .Generate(Generate[9]) );
  PG_generate_7 PG_GEN_10__PG_generate_inst ( .add_1(add_1[10]), .add_2(
        add_2[10]), .Propagate(Propagate[10]), .Generate(Generate[10]) );
  PG_generate_6 PG_GEN_11__PG_generate_inst ( .add_1(add_1[11]), .add_2(
        add_2[11]), .Propagate(Propagate[11]), .Generate(Generate[11]) );
  PG_generate_5 PG_GEN_12__PG_generate_inst ( .add_1(add_1[12]), .add_2(
        add_2[12]), .Propagate(Propagate[12]), .Generate(Generate[12]) );
  PG_generate_4 PG_GEN_13__PG_generate_inst ( .add_1(add_1[13]), .add_2(
        add_2[13]), .Propagate(Propagate[13]), .Generate(Generate[13]) );
  PG_generate_3 PG_GEN_14__PG_generate_inst ( .add_1(add_1[14]), .add_2(
        add_2[14]), .Propagate(Propagate[14]), .Generate(Generate[14]) );
  PG_generate_2 PG_GEN_15__PG_generate_inst ( .add_1(add_1[15]), .add_2(
        add_2[15]), .Propagate(Propagate[15]), .Generate(Generate[15]) );
  PG_generate_1 PG_GEN_16__PG_generate_inst ( .add_1(add_1[16]), .add_2(
        add_2[16]), .Propagate(Propagate[16]), .Generate(Generate[16]) );
  CUS_PLUS_0 STAGE_1_GEN_2__STAGE_1_GEN_CUS_PLUS_inst ( .g_high(Generate[2]), 
        .g_low(Generate[1]), .p_high(Propagate[2]), .p_low(Propagate[1]), 
        .alpha(stage_1_alpha_2), .beta(stage_1_beta_2) );
  CUS_PLUS_25 STAGE_1_GEN_4__STAGE_1_GEN_CUS_PLUS_inst ( .g_high(Generate[4]), 
        .g_low(Generate[3]), .p_high(Propagate[4]), .p_low(Propagate[3]), 
        .alpha(stage_1_alpha_4), .beta(stage_1_beta_4) );
  CUS_PLUS_24 STAGE_1_GEN_6__STAGE_1_GEN_CUS_PLUS_inst ( .g_high(Generate[6]), 
        .g_low(Generate[5]), .p_high(Propagate[6]), .p_low(Propagate[5]), 
        .alpha(stage_1_alpha_6), .beta(stage_1_beta_6) );
  CUS_PLUS_23 STAGE_1_GEN_8__STAGE_1_GEN_CUS_PLUS_inst ( .g_high(Generate[8]), 
        .g_low(Generate[7]), .p_high(Propagate[8]), .p_low(Propagate[7]), 
        .alpha(stage_1_alpha_8), .beta(stage_1_beta_8) );
  CUS_PLUS_22 STAGE_1_GEN_10__STAGE_1_GEN_CUS_PLUS_inst ( .g_high(Generate[10]), .g_low(Generate[9]), .p_high(Propagate[10]), .p_low(Propagate[9]), .alpha(
        stage_1_alpha_10), .beta(stage_1_beta_10) );
  CUS_PLUS_21 STAGE_1_GEN_12__STAGE_1_GEN_CUS_PLUS_inst ( .g_high(Generate[12]), .g_low(Generate[11]), .p_high(Propagate[12]), .p_low(Propagate[11]), .alpha(
        stage_1_alpha_12), .beta(stage_1_beta_12) );
  CUS_PLUS_20 STAGE_1_GEN_14__STAGE_1_GEN_CUS_PLUS_inst ( .g_high(Generate[14]), .g_low(Generate[13]), .p_high(Propagate[14]), .p_low(Propagate[13]), .alpha(
        stage_1_alpha_14), .beta(stage_1_beta_14) );
  CUS_PLUS_19 STAGE_1_GEN_16__STAGE_1_GEN_CUS_PLUS_inst ( .g_high(Generate[16]), .g_low(Generate[15]), .p_high(Propagate[16]), .p_low(Propagate[15]), .alpha(
        stage_1_alpha_16_), .beta(stage_1_beta_16_) );
  CUS_PLUS_18 STAGE_2_GEN_4__STAGE_2_GEN_CUS_PLUS_inst ( .g_high(
        stage_1_alpha_4), .g_low(stage_1_alpha_2), .p_high(stage_1_beta_4), 
        .p_low(stage_1_beta_2), .alpha(stage_2_alpha_4), .beta(stage_2_beta_4)
         );
  CUS_PLUS_17 STAGE_2_GEN_8__STAGE_2_GEN_CUS_PLUS_inst ( .g_high(
        stage_1_alpha_8), .g_low(stage_1_alpha_6), .p_high(stage_1_beta_8), 
        .p_low(stage_1_beta_6), .alpha(stage_2_alpha_8), .beta(stage_2_beta_8)
         );
  CUS_PLUS_16 STAGE_2_GEN_12__STAGE_2_GEN_CUS_PLUS_inst ( .g_high(
        stage_1_alpha_12), .g_low(stage_1_alpha_10), .p_high(stage_1_beta_12), 
        .p_low(stage_1_beta_10), .alpha(stage_2_alpha_12), .beta(
        stage_2_beta_12) );
  CUS_PLUS_15 STAGE_2_GEN_16__STAGE_2_GEN_CUS_PLUS_inst ( .g_high(
        stage_1_alpha_16_), .g_low(stage_1_alpha_14), .p_high(stage_1_beta_16_), .p_low(stage_1_beta_14), .alpha(stage_2_alpha_16_), .beta(stage_2_beta_16_)
         );
  CUS_PLUS_14 STAGE_3_GEN_8__STAGE_3_GEN_CUS_PLUS_inst ( .g_high(
        stage_2_alpha_8), .g_low(stage_2_alpha_4), .p_high(stage_2_beta_8), 
        .p_low(stage_2_beta_4), .alpha(stage_3_alpha_8), .beta(stage_3_beta_8)
         );
  CUS_PLUS_13 STAGE_3_GEN_16__STAGE_3_GEN_CUS_PLUS_inst ( .g_high(
        stage_2_alpha_16_), .g_low(stage_2_alpha_12), .p_high(stage_2_beta_16_), .p_low(stage_2_beta_12), .alpha(stage_3_alpha_16_), .beta(stage_3_beta_16_)
         );
  CUS_PLUS_12 STAGE_4_GEN_12__STAGE_4_GEN_CUS_PLUS_inst ( .g_high(
        stage_2_alpha_12), .g_low(stage_3_alpha_8), .p_high(stage_2_beta_12), 
        .p_low(stage_3_beta_8), .alpha(stage_4_alpha_12), .beta(
        stage_4_beta_12) );
  CUS_PLUS_11 STAGE_4_GEN_16__STAGE_4_GEN_CUS_PLUS_inst ( .g_high(
        stage_3_alpha_16_), .g_low(stage_3_alpha_8), .p_high(stage_3_beta_16_), 
        .p_low(stage_3_beta_8), .alpha(stage_4_alpha_16_), .beta(
        stage_4_beta_16_) );
  CUS_PLUS_10 STAGE_5_GEN_6__STAGE_5_GEN_CUS_PLUS_inst ( .g_high(
        stage_1_alpha_6), .g_low(stage_2_alpha_4), .p_high(stage_1_beta_6), 
        .p_low(stage_2_beta_4), .alpha(stage_5_alpha_6), .beta(stage_5_beta_6)
         );
  CUS_PLUS_9 STAGE_5_GEN_10__STAGE_5_GEN_CUS_PLUS_inst ( .g_high(
        stage_1_alpha_10), .g_low(stage_3_alpha_8), .p_high(stage_1_beta_10), 
        .p_low(stage_3_beta_8), .alpha(stage_5_alpha_10), .beta(
        stage_5_beta_10) );
  CUS_PLUS_8 STAGE_5_GEN_14__STAGE_5_GEN_CUS_PLUS_inst ( .g_high(
        stage_1_alpha_14), .g_low(stage_4_alpha_12), .p_high(stage_1_beta_14), 
        .p_low(stage_4_beta_12), .alpha(stage_5_alpha_14_), .beta(
        stage_5_beta_14_) );
  CUS_PLUS_7 STAGE_6_GEN_3__STAGE_6_GEN_CUS_PLUS_inst ( .g_high(Generate[3]), 
        .g_low(stage_1_alpha_2), .p_high(Propagate[3]), .p_low(stage_1_beta_2), 
        .alpha(stage_6_alpha_3), .beta(stage_6_beta_3) );
  CUS_PLUS_6 STAGE_6_GEN_5__STAGE_6_GEN_CUS_PLUS_inst ( .g_high(Generate[5]), 
        .g_low(stage_2_alpha_4), .p_high(Propagate[5]), .p_low(stage_2_beta_4), 
        .alpha(stage_6_alpha_5), .beta(stage_6_beta_5) );
  CUS_PLUS_5 STAGE_6_GEN_7__STAGE_6_GEN_CUS_PLUS_inst ( .g_high(Generate[7]), 
        .g_low(stage_5_alpha_6), .p_high(Propagate[7]), .p_low(stage_5_beta_6), 
        .alpha(stage_6_alpha_7), .beta(stage_6_beta_7) );
  CUS_PLUS_4 STAGE_6_GEN_9__STAGE_6_GEN_CUS_PLUS_inst ( .g_high(Generate[9]), 
        .g_low(stage_3_alpha_8), .p_high(Propagate[9]), .p_low(stage_3_beta_8), 
        .alpha(stage_6_alpha_9), .beta(stage_6_beta_9) );
  CUS_PLUS_3 STAGE_6_GEN_11__STAGE_6_GEN_CUS_PLUS_inst ( .g_high(Generate[11]), 
        .g_low(stage_5_alpha_10), .p_high(Propagate[11]), .p_low(
        stage_5_beta_10), .alpha(stage_6_alpha_11), .beta(stage_6_beta_11) );
  CUS_PLUS_2 STAGE_6_GEN_13__STAGE_6_GEN_CUS_PLUS_inst ( .g_high(Generate[13]), 
        .g_low(stage_4_alpha_12), .p_high(Propagate[13]), .p_low(
        stage_4_beta_12), .alpha(stage_6_alpha_13), .beta(stage_6_beta_13) );
  CUS_PLUS_1 STAGE_6_GEN_15__STAGE_6_GEN_CUS_PLUS_inst ( .g_high(Generate[15]), 
        .g_low(stage_5_alpha_14_), .p_high(Propagate[15]), .p_low(
        stage_5_beta_14_), .alpha(stage_6_alpha_15_), .beta(stage_6_beta_15_)
         );
  Carry_Generate_0 CARRY_GEN_1__Carry_Generate_inst ( .alpha(Generate[1]), 
        .beta(Propagate[1]), .c_in(c_in), .c_out(Carry[1]) );
  Carry_Generate_15 CARRY_GEN_2__Carry_Generate_inst ( .alpha(stage_1_alpha_2), 
        .beta(stage_1_beta_2), .c_in(Carry[1]), .c_out(Carry[2]) );
  Carry_Generate_14 CARRY_GEN_3__Carry_Generate_inst ( .alpha(stage_6_alpha_3), 
        .beta(stage_6_beta_3), .c_in(Carry[2]), .c_out(Carry[3]) );
  Carry_Generate_13 CARRY_GEN_4__Carry_Generate_inst ( .alpha(stage_2_alpha_4), 
        .beta(stage_2_beta_4), .c_in(Carry[3]), .c_out(Carry[4]) );
  Carry_Generate_12 CARRY_GEN_5__Carry_Generate_inst ( .alpha(stage_6_alpha_5), 
        .beta(stage_6_beta_5), .c_in(Carry[4]), .c_out(Carry[5]) );
  Carry_Generate_11 CARRY_GEN_6__Carry_Generate_inst ( .alpha(stage_5_alpha_6), 
        .beta(stage_5_beta_6), .c_in(Carry[5]), .c_out(Carry[6]) );
  Carry_Generate_10 CARRY_GEN_7__Carry_Generate_inst ( .alpha(stage_6_alpha_7), 
        .beta(stage_6_beta_7), .c_in(Carry[6]), .c_out(Carry[7]) );
  Carry_Generate_9 CARRY_GEN_8__Carry_Generate_inst ( .alpha(stage_3_alpha_8), 
        .beta(stage_3_beta_8), .c_in(Carry[7]), .c_out(Carry[8]) );
  Carry_Generate_8 CARRY_GEN_9__Carry_Generate_inst ( .alpha(stage_6_alpha_9), 
        .beta(stage_6_beta_9), .c_in(Carry[8]), .c_out(Carry[9]) );
  Carry_Generate_7 CARRY_GEN_10__Carry_Generate_inst ( .alpha(stage_5_alpha_10), .beta(stage_5_beta_10), .c_in(Carry[9]), .c_out(Carry[10]) );
  Carry_Generate_6 CARRY_GEN_11__Carry_Generate_inst ( .alpha(stage_6_alpha_11), .beta(stage_6_beta_11), .c_in(Carry[10]), .c_out(Carry[11]) );
  Carry_Generate_5 CARRY_GEN_12__Carry_Generate_inst ( .alpha(stage_4_alpha_12), .beta(stage_4_beta_12), .c_in(Carry[11]), .c_out(Carry[12]) );
  Carry_Generate_4 CARRY_GEN_13__Carry_Generate_inst ( .alpha(stage_6_alpha_13), .beta(stage_6_beta_13), .c_in(Carry[12]), .c_out(Carry[13]) );
  Carry_Generate_3 CARRY_GEN_14__Carry_Generate_inst ( .alpha(
        stage_5_alpha_14_), .beta(stage_5_beta_14_), .c_in(Carry[13]), .c_out(
        Carry[14]) );
  Carry_Generate_2 CARRY_GEN_15__Carry_Generate_inst ( .alpha(
        stage_6_alpha_15_), .beta(stage_6_beta_15_), .c_in(Carry[14]), .c_out(
        Carry[15]) );
  Carry_Generate_1 CARRY_GEN_16__Carry_Generate_inst ( .alpha(
        stage_4_alpha_16_), .beta(stage_4_beta_16_), .c_in(Carry[15]), .c_out(
        c_out[0]) );
  SUM_generate_0 SUM_GEN_1__SUM_generate_inst ( .Propagate(Propagate[1]), 
        .c_in(c_in), .Sum(sum[1]) );
  SUM_generate_15 SUM_GEN_2__SUM_generate_inst ( .Propagate(Propagate[2]), 
        .c_in(Carry[1]), .Sum(sum[2]) );
  SUM_generate_14 SUM_GEN_3__SUM_generate_inst ( .Propagate(Propagate[3]), 
        .c_in(Carry[2]), .Sum(sum[3]) );
  SUM_generate_13 SUM_GEN_4__SUM_generate_inst ( .Propagate(Propagate[4]), 
        .c_in(Carry[3]), .Sum(sum[4]) );
  SUM_generate_12 SUM_GEN_5__SUM_generate_inst ( .Propagate(Propagate[5]), 
        .c_in(Carry[4]), .Sum(sum[5]) );
  SUM_generate_11 SUM_GEN_6__SUM_generate_inst ( .Propagate(Propagate[6]), 
        .c_in(Carry[5]), .Sum(sum[6]) );
  SUM_generate_10 SUM_GEN_7__SUM_generate_inst ( .Propagate(Propagate[7]), 
        .c_in(Carry[6]), .Sum(sum[7]) );
  SUM_generate_9 SUM_GEN_8__SUM_generate_inst ( .Propagate(Propagate[8]), 
        .c_in(Carry[7]), .Sum(sum[8]) );
  SUM_generate_8 SUM_GEN_9__SUM_generate_inst ( .Propagate(Propagate[9]), 
        .c_in(Carry[8]), .Sum(sum[9]) );
  SUM_generate_7 SUM_GEN_10__SUM_generate_inst ( .Propagate(Propagate[10]), 
        .c_in(Carry[9]), .Sum(sum[10]) );
  SUM_generate_6 SUM_GEN_11__SUM_generate_inst ( .Propagate(Propagate[11]), 
        .c_in(Carry[10]), .Sum(sum[11]) );
  SUM_generate_5 SUM_GEN_12__SUM_generate_inst ( .Propagate(Propagate[12]), 
        .c_in(Carry[11]), .Sum(sum[12]) );
  SUM_generate_4 SUM_GEN_13__SUM_generate_inst ( .Propagate(Propagate[13]), 
        .c_in(Carry[12]), .Sum(sum[13]) );
  SUM_generate_3 SUM_GEN_14__SUM_generate_inst ( .Propagate(Propagate[14]), 
        .c_in(Carry[13]), .Sum(sum[14]) );
  SUM_generate_2 SUM_GEN_15__SUM_generate_inst ( .Propagate(Propagate[15]), 
        .c_in(Carry[14]), .Sum(sum[15]) );
  SUM_generate_1 SUM_GEN_16__SUM_generate_inst ( .Propagate(Propagate[16]), 
        .c_in(Carry[15]), .Sum(sum[16]) );
endmodule

