module one_bit_full_adder
